module memory(A, B)