module controller(clk, rst);
    input wire clk, rst;

    
endmodule